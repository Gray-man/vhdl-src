library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_signed.all;
use IEEE.numeric_std.all;

entity data_path is
port(
	    );
end entity data_path;

architecture data_path of data_path is

begin
	regfile: entity work.regfile




end architecture data_path;
















